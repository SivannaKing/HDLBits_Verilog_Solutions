module top_module (
    input clk,
    input [7:0] in,
    output [7:0] pedge
);

	reg [7:0] d_last;	
	// TODO IMP posedge detect
	always @(posedge clk) begin
		d_last <= in;			// Remember the state of the previous cycle
		pedge <= in & ~d_last;	// A positive edge occurred if input was 0 and is now 1.
	end
    
endmodule