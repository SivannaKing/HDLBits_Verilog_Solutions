// Note the Verilog-1995 module declaration syntax here:
module top_module (
    clk,
    reset,
    in,
    out
);
    input clk;
    input reset;  // Synchronous reset to state B
    input in;
    output out;  //  
    reg out;

    // Fill in state name declarations
    parameter A = 0, B = 1;
    reg present_state, next_state;
    //组合电路
    always @(*) begin
        case (present_state)
            // Fill in state transition logic
            A: next_state = in ? A : B;
            B: next_state = in ? B : A;
        endcase
    end
    //时序电路
    always @(posedge clk) begin
        if (reset) begin
            // Fill in reset logic
            present_state <= B;
        end else present_state <= next_state;
    end
    assign out = present_state;
endmodule
